// -- python C:\Users\Brandon\Documents\Personal_Projects\my_utils\modelsim_utils\auto_run.py -d run_cmd__nand4_gate_v.do

module not1_gate_v
  (input i_a,
   output o_f);
   
  assign o_f = ~i_a;
  
endmodule







